module adder32(op1, op2, control, Output);
	input [31:0] op1, op2;
	input control;
	output [31:0] Output;
	
	
endmodule 